`timescale 1ns / 1ps

module TLlab6(

    );
    
    
endmodule

